`timescale 1ns / 1ps
//Source: http://www.bigmessowires.com/2009/06/21/fpga-pong/
//modified to run on the new CRT driver
//and 100MHz system clock
//ECE433 Fall 2022
// -----------------------------------------------
// updates the ball and paddle positions, and
// determines the output video image
// -----------------------------------------------
module game2022fallTemplate(
input Reset, clk25, rota, rotb,
input [9:0] xpos, ypos,
output [3:0] red, green, blue);
		
		
endmodule
